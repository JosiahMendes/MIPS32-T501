module test();
endmodule