module cpu_bus_tb;
    logic clock;
    logic rst;


endmodule