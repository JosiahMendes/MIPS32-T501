module cpu_bus_tb.v;
    logic clock;
    logic reset;



endmodule
